`timescale 1ns / 1ps

module tb();
  always // always_comb, always_ff, always_latch
    always statement;
  always begin
  ...
  end
  
endmodule