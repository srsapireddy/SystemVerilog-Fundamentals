// Create Monitor and Scoreboard Code for Synchronous 4-bit Multiplier. Stimulus is generated in Testbench top so do not add Transaction, 
// Generator, or Driver Code. Also, add the Scoreboard model to compare the response with an expected result.
