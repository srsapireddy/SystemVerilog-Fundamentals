class first;
  bit [2:0] data;
  bit [1:0] data2;
  
endclass

module tb;
  first f;
  f.data;
  f.data2;
endmodule